`timescale 1ns/100ps

module Compare (A, B, Y);

endmodule
